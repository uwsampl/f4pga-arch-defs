`default_nettype none
module PUR(input PUR);
    parameter RST_PULSE;
endmodule
