`default_nettype none
module GSR(input GSR);
endmodule
