`default_nettype none
module IB(input I, output O);
    assign O = I;
endmodule
