`default_nettype none
module OB(input I, output O);
    assign O = I;
endmodule
